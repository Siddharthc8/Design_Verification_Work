package axi_env_pkg;


import uvm_pkg::*;

`include "transaction.sv"
`include "reset_sequence.sv"
`include "incr_sequence.sv"
`include "fixed_sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "imonitor.sv"
`include "master_agent.sv"
`include "omonitor.sv"
`include "slave_agent.sv"
`include "scoreboard.sv"
`include "environment.sv"

endpackage
